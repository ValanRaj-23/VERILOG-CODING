module top_module ( input x, input y, output z );
    
    xnor G0(z, x, y);

endmodule
